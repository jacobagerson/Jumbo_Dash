--library IEEE;
--use IEEE.std_logic_1164.all;
--use IEEE.numeric_std.all;


--entity ground3ROM is
--port(
	--Xin : in unsigned(4 downto 0);
	--Yin : in unsigned(4 downto 0);
--data : out std_logic_vector(5 downto 0)
--);
--end entity;


--architecture synth of ground3ROM is


--Signal addy : unsigned(9 downto 0);


--Begin


--addy <= Yin & Xin;


--process(addy) begin
	--case addy is
		--when "0000101101" => data <= "000000";
--when "0000101110" => data <= "000000";
--when "0000101111" => data <= "000000";
--when "0000110000" => data <= "000000";
--when "0000110001" => data <= "000000";
--when "0000110010" => data <= "000000";
--when "0000110011" => data <= "000000";
--when "0000110100" => data <= "000000";
--when "0000110101" => data <= "000000";
--when "0001001011" => data <= "000000";
--when "0001001100" => data <= "000000";
--when "0001001101" => data <= "000000";
--when "0001010101" => data <= "000000";
--when "0001010110" => data <= "000000";
--when "0001100000" => data <= "000000";
--when "0001100001" => data <= "000000";
--when "0001100010" => data <= "000000";
--when "0001100011" => data <= "000000";
--when "0001100100" => data <= "000000";
--when "0001100101" => data <= "000000";
--when "0001100110" => data <= "000000";
--when "0001100111" => data <= "000000";
--when "0001101000" => data <= "000000";
--when "0001101001" => data <= "000000";
--when "0001101010" => data <= "000000";
--when "0001101011" => data <= "000000";
--when "0001110110" => data <= "000000";
--when "0001110111" => data <= "000000";
--when "0001111000" => data <= "000000";
--when "0001111001" => data <= "000000";
--when "0001111010" => data <= "000000";
--when "0001111011" => data <= "000000";
--when "0001111100" => data <= "000000";
--when "0001111101" => data <= "000000";
--when "0001111110" => data <= "000000";
--when "0011010000" => data <= "000000";
--when "0011100101" => data <= "000000";
--when "0011100110" => data <= "000000";
--when "0011100111" => data <= "000000";
--when "0011101000" => data <= "000000";
--when "0100011000" => data <= "000000";
--when "0100011001" => data <= "000000";
--when "0101001100" => data <= "000000";
--when "0110010111" => data <= "000000";
--when "0110011000" => data <= "000000";
--when "0110100011" => data <= "000000";
		--when others => data <= "111111";
--end case;
--end process;
--end;











