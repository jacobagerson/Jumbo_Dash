--library IEEE;
--use IEEE.std_logic_1164.all;
--use IEEE.numeric_std.all;


--entity ground4ROM is
--port(
	--Xin : in unsigned(4 downto 0);
	--Yin : in unsigned(4 downto 0);
--data : out std_logic_vector(5 downto 0)
--);
--end entity;


--architecture synth of ground4ROM is


--Signal addy : unsigned(9 downto 0);


--Begin


--addy <= Yin & Xin;


--process(addy) begin
	--case addy is
		--when "0000110110" => data <= "000000";
--when "0000110111" => data <= "000000";
--when "0000111000" => data <= "000000";
--when "0000111001" => data <= "000000";
--when "0001010100" => data <= "000000";
--when "0001010101" => data <= "000000";
--when "0001010110" => data <= "000000";
--when "0001011001" => data <= "000000";
--when "0001011010" => data <= "000000";
--when "0001011011" => data <= "000000";
--when "0001100000" => data <= "000000";
--when "0001100001" => data <= "000000";
--when "0001100010" => data <= "000000";
--when "0001100011" => data <= "000000";
--when "0001110011" => data <= "000000";
--when "0001110100" => data <= "000000";
--when "0001111011" => data <= "000000";
--when "0001111100" => data <= "000000";
--when "0001111101" => data <= "000000";
--when "0001111110" => data <= "000000";
--when "0010000011" => data <= "000000";
--when "0010000100" => data <= "000000";
--when "0010000101" => data <= "000000";
--when "0010000110" => data <= "000000";
--when "0010000111" => data <= "000000";
--when "0010001000" => data <= "000000";
--when "0010001101" => data <= "000000";
--when "0010001110" => data <= "000000";
--when "0010001111" => data <= "000000";
--when "0010010000" => data <= "000000";
--when "0010010001" => data <= "000000";
--when "0010010010" => data <= "000000";
--when "0010010011" => data <= "000000";
--when "0010101000" => data <= "000000";
--when "0010101001" => data <= "000000";
--when "0010101010" => data <= "000000";
--when "0010101011" => data <= "000000";
--when "0010101100" => data <= "000000";
--when "0010101101" => data <= "000000";
--when "0011110111" => data <= "000000";
--when "0011111000" => data <= "000000";
--when "0100000010" => data <= "000000";
--when "0100000011" => data <= "000000";
--when "0100110001" => data <= "000000";
--when "0101101000" => data <= "000000";
--when "0101101001" => data <= "000000";
--when "0101101010" => data <= "000000";
--when "0101111010" => data <= "000000";
--when "0111010100" => data <= "000000";
--when "0111010101" => data <= "000000";
		--when others => data <= "111111";
--end case;
--end process;
--end;











