library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity pterodown_ROM is
port(
	Xin : in unsigned(4 downto 0);
	Yin : in unsigned(4 downto 0);
data : out std_logic_vector(5 downto 0)
);
end pterodown_ROM;


architecture synth of pterodown_ROM is

signal addy : unsigned(9 downto 0);
begin

addy <= Yin & Xin;

process(addy) begin
	case addy is
		when "0010100100" => data <= "000000";
when "0010100101" => data <= "000000";
when "0011000011" => data <= "000000";
when "0011000100" => data <= "000000";
when "0011000101" => data <= "000000";
when "0011000110" => data <= "000000";
when "0011100010" => data <= "000000";
when "0011100011" => data <= "000000";
when "0011100100" => data <= "000000";
when "0011100101" => data <= "000000";
when "0011100110" => data <= "000000";
when "0011100111" => data <= "000000";
when "0100000001" => data <= "000000";
when "0100000010" => data <= "000000";
when "0100000011" => data <= "000000";
when "0100000100" => data <= "000000";
when "0100000101" => data <= "000000";
when "0100000110" => data <= "000000";
when "0100000111" => data <= "000000";
when "0100100000" => data <= "000000";
when "0100100001" => data <= "000000";
when "0100100010" => data <= "000000";
when "0100100011" => data <= "000000";
when "0100100100" => data <= "000000";
when "0100100101" => data <= "000000";
when "0100100110" => data <= "000000";
when "0100100111" => data <= "000000";
when "0100101000" => data <= "000000";
when "0100101001" => data <= "000000";
when "0100101010" => data <= "000000";
when "0100101011" => data <= "000000";
when "0100101100" => data <= "000000";
when "0100101101" => data <= "000000";
when "0100101110" => data <= "000000";
when "0100101111" => data <= "000000";
when "0100110000" => data <= "000000";
when "0100110001" => data <= "000000";
when "0100110010" => data <= "000000";
when "0100110011" => data <= "000000";
when "0100110100" => data <= "000000";
when "0101000101" => data <= "000000";
when "0101000110" => data <= "000000";
when "0101000111" => data <= "000000";
when "0101001000" => data <= "000000";
when "0101001001" => data <= "000000";
when "0101001010" => data <= "000000";
when "0101001011" => data <= "000000";
when "0101001100" => data <= "000000";
when "0101001101" => data <= "000000";
when "0101001110" => data <= "000000";
when "0101001111" => data <= "000000";
when "0101010000" => data <= "000000";
when "0101010001" => data <= "000000";
when "0101100111" => data <= "000000";
when "0101101000" => data <= "000000";
when "0101101001" => data <= "000000";
when "0101101010" => data <= "000000";
when "0101101011" => data <= "000000";
when "0101101100" => data <= "000000";
when "0101101101" => data <= "000000";
when "0101101110" => data <= "000000";
when "0101101111" => data <= "000000";
when "0101110000" => data <= "000000";
when "0101110001" => data <= "000000";
when "0101110010" => data <= "000000";
when "0101110011" => data <= "000000";
when "0110001001" => data <= "000000";
when "0110001010" => data <= "000000";
when "0110001011" => data <= "000000";
when "0110001100" => data <= "000000";
when "0110001101" => data <= "000000";
when "0110001110" => data <= "000000";
when "0110001111" => data <= "000000";
when "0110010000" => data <= "000000";
when "0110101001" => data <= "000000";
when "0110101010" => data <= "000000";
when "0110101011" => data <= "000000";
when "0110101100" => data <= "000000";
when "0110101101" => data <= "000000";
when "0110101110" => data <= "000000";
when "0110101111" => data <= "000000";
when "0111001001" => data <= "000000";
when "0111001010" => data <= "000000";
when "0111001011" => data <= "000000";
when "0111001100" => data <= "000000";
when "0111001101" => data <= "000000";
when "0111001110" => data <= "000000";
when "0111101001" => data <= "000000";
when "0111101010" => data <= "000000";
when "0111101011" => data <= "000000";
when "0111101100" => data <= "000000";
when "0111101101" => data <= "000000";
when "1000001001" => data <= "000000";
when "1000001010" => data <= "000000";
when "1000001011" => data <= "000000";
when "1000001100" => data <= "000000";
when "1000101001" => data <= "000000";
when "1000101010" => data <= "000000";
when "1000101011" => data <= "000000";
when "1001001001" => data <= "000000";
when "1001001010" => data <= "000000";
when "1001101001" => data <= "000000";
when others => data <= "111111";


end case;
end process;
end;
