--library IEEE;
--use IEEE.std_logic_1164.all;
--use IEEE.numeric_std.all;


--entity ground2ROM is
--port(
	--Xin : in unsigned(4 downto 0);
	--Yin : in unsigned(4 downto 0);
--data : out std_logic_vector(5 downto 0)
--);
--end entity;


--architecture synth of ground2ROM is


--Signal addy : unsigned(9 downto 0);


--Begin


--addy <= Yin & Xin;


--process(addy) begin
	--case addy is
		--when "0001010001" => data <= "000000";
--when "0001010010" => data <= "000000";
--when "0001010011" => data <= "000000";
--when "0001010100" => data <= "000000";
--when "0001010101" => data <= "000000";
--when "0001010110" => data <= "000000";
--when "0001100000" => data <= "000000";
--when "0001100001" => data <= "000000";
--when "0001100010" => data <= "000000";
--when "0001100011" => data <= "000000";
--when "0001100100" => data <= "000000";
--when "0001100101" => data <= "000000";
--when "0001101100" => data <= "000000";
--when "0001101101" => data <= "000000";
--when "0001101110" => data <= "000000";
--when "0001101111" => data <= "000000";
--when "0001110000" => data <= "000000";
--when "0001110001" => data <= "000000";
--when "0001110110" => data <= "000000";
--when "0001110111" => data <= "000000";
--when "0001111000" => data <= "000000";
--when "0001111011" => data <= "000000";
--when "0001111100" => data <= "000000";
--when "0001111101" => data <= "000000";
--when "0001111110" => data <= "000000";
--when "0010000101" => data <= "000000";
--when "0010000110" => data <= "000000";
--when "0010001011" => data <= "000000";
--when "0010001100" => data <= "000000";
--when "0010011000" => data <= "000000";
--when "0010011001" => data <= "000000";
--when "0010011010" => data <= "000000";
--when "0010011011" => data <= "000000";
--when "0010100110" => data <= "000000";
--when "0010100111" => data <= "000000";
--when "0010101000" => data <= "000000";
--when "0010101001" => data <= "000000";
--when "0010101010" => data <= "000000";
--when "0010101011" => data <= "000000";
--when "0011111011" => data <= "000000";
--when "0100110010" => data <= "000000";
--when "0100110011" => data <= "000000";
--when "0100110100" => data <= "000000";
--when "0101000011" => data <= "000000";
--when "0101000100" => data <= "000000";
--when "0101000101" => data <= "000000";
--when "0110011011" => data <= "000000";
--when "0110101110" => data <= "000000";
		--when others => data <= "111111";
--end case;
--end process;
--end;











