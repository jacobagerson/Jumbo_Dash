library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity CactusROM4 is
	port(
		Xin : in unsigned(4 downto 0);
		Yin : in unsigned(4 downto 0);
		data : out std_logic_vector(5 downto 0)
	);
end CactusROM4;

architecture synth of CactusROM4 is
	signal addy : unsigned(9 downto 0);

begin
	addy <= Yin & Xin;

	process(addy) begin
		case addy is
			when "0000000100" => data <= "000000";
			when "0000100011" => data <= "000000";
			when "0000100100" => data <= "000000";
			when "0000100101" => data <= "000000";
			when "0001000011" => data <= "000000";
			when "0001000100" => data <= "000000";
			when "0001000101" => data <= "000000";
			when "0001001000" => data <= "000000";
			when "0001100011" => data <= "000000";
			when "0001100100" => data <= "000000";
			when "0001100101" => data <= "000000";
			when "0001100111" => data <= "000000";
			when "0001101000" => data <= "000000";
			when "0010000001" => data <= "000000";
			when "0010000011" => data <= "000000";
			when "0010000100" => data <= "000000";
			when "0010000101" => data <= "000000";
			when "0010000111" => data <= "000000";
			when "0010001000" => data <= "000000";
			when "0010100000" => data <= "000000";
			when "0010100001" => data <= "000000";
			when "0010100011" => data <= "000000";
			when "0010100100" => data <= "000000";
			when "0010100101" => data <= "000000";
			when "0010100111" => data <= "000000";
			when "0010101000" => data <= "000000";
			when "0011000000" => data <= "000000";
			when "0011000001" => data <= "000000";
			when "0011000011" => data <= "000000";
			when "0011000100" => data <= "000000";
			when "0011000101" => data <= "000000";
			when "0011000111" => data <= "000000";
			when "0011001000" => data <= "000000";
			when "0011100000" => data <= "000000";
			when "0011100001" => data <= "000000";
			when "0011100011" => data <= "000000";
			when "0011100100" => data <= "000000";
			when "0011100101" => data <= "000000";
			when "0011100111" => data <= "000000";
			when "0011101000" => data <= "000000";
			when "0100000000" => data <= "000000";
			when "0100000001" => data <= "000000";
			when "0100000011" => data <= "000000";
			when "0100000100" => data <= "000000";
			when "0100000101" => data <= "000000";
			when "0100000110" => data <= "000000";
			when "0100000111" => data <= "000000";
			when "0100001000" => data <= "000000";
			when "0100100000" => data <= "000000";
			when "0100100001" => data <= "000000";
			when "0100100011" => data <= "000000";
			when "0100100100" => data <= "000000";
			when "0100100101" => data <= "000000";
			when "0100100110" => data <= "000000";
			when "0100100111" => data <= "000000";
			when "0101000000" => data <= "000000";
			when "0101000001" => data <= "000000";
			when "0101000011" => data <= "000000";
			when "0101000100" => data <= "000000";
			when "0101000101" => data <= "000000";
			when "0101100000" => data <= "000000";
			when "0101100001" => data <= "000000";
			when "0101100011" => data <= "000000";
			when "0101100100" => data <= "000000";
			when "0101100101" => data <= "000000";
			when "0110000000" => data <= "000000";
			when "0110000001" => data <= "000000";
			when "0110000011" => data <= "000000";
			when "0110000100" => data <= "000000";
			when "0110000101" => data <= "000000";
			when "0110100000" => data <= "000000";
			when "0110100001" => data <= "000000";
			when "0110100011" => data <= "000000";
			when "0110100100" => data <= "000000";
			when "0110100101" => data <= "000000";
			when "0111000000" => data <= "000000";
			when "0111000001" => data <= "000000";
			when "0111000010" => data <= "000000";
			when "0111000011" => data <= "000000";
			when "0111000100" => data <= "000000";
			when "0111000101" => data <= "000000";
			when "0111100001" => data <= "000000";
			when "0111100010" => data <= "000000";
			when "0111100011" => data <= "000000";
			when "0111100100" => data <= "000000";
			when "0111100101" => data <= "000000";
			when "1000000011" => data <= "000000";
			when "1000000100" => data <= "000000";
			when "1000000101" => data <= "000000";
			when "1000100011" => data <= "000000";
			when "1000100100" => data <= "000000";
			when "1000100101" => data <= "000000";
			when "1001000011" => data <= "000000";
			when "1001000100" => data <= "000000";
			when "1001000101" => data <= "000000";
			when "1001100011" => data <= "000000";
			when "1001100100" => data <= "000000";
			when "1001100101" => data <= "000000";
			when "1010000011" => data <= "000000";
			when "1010000100" => data <= "000000";
			when "1010000101" => data <= "000000";
			when others => data <= "111111";
		end case;
	end process;
end synth;
