--library IEEE;
--use IEEE.std_logic_1164.all;
--use IEEE.numeric_std.all;


--entity ground5ROM is
--port(
	--Xin : in unsigned(4 downto 0);
	--Yin : in unsigned(4 downto 0);
--data : out std_logic_vector(5 downto 0)
--);
--end entity;


--architecture synth of ground5ROM is


--Signal addy : unsigned(9 downto 0);


--Begin


--addy <= Yin & Xin;


--process(addy) begin
	--case addy is
		--when "0001100000" => data <= "000000";
--when "0001100001" => data <= "000000";
--when "0001100010" => data <= "000000";
--when "0001100011" => data <= "000000";
--when "0001100100" => data <= "000000";
--when "0001100101" => data <= "000000";
--when "0001100110" => data <= "000000";
--when "0001100111" => data <= "000000";
--when "0001110011" => data <= "000000";
--when "0001110100" => data <= "000000";
--when "0001110101" => data <= "000000";
--when "0001110110" => data <= "000000";
--when "0001110111" => data <= "000000";
--when "0001111000" => data <= "000000";
--when "0001111001" => data <= "000000";
--when "0001111010" => data <= "000000";
--when "0001111011" => data <= "000000";
--when "0001111100" => data <= "000000";
--when "0001111101" => data <= "000000";
--when "0001111110" => data <= "000000";
--when "0010000111" => data <= "000000";
--when "0010001000" => data <= "000000";
--when "0010001001" => data <= "000000";
--when "0010001010" => data <= "000000";
--when "0010001111" => data <= "000000";
--when "0010010000" => data <= "000000";
--when "0010010001" => data <= "000000";
--when "0010010010" => data <= "000000";
--when "0010010011" => data <= "000000";
--when "0010101010" => data <= "000000";
--when "0010101011" => data <= "000000";
--when "0010101100" => data <= "000000";
--when "0010101101" => data <= "000000";
--when "0010101110" => data <= "000000";
--when "0010101111" => data <= "000000";
--when "0011110011" => data <= "000000";
--when "0100000110" => data <= "000000";
--when "0100000111" => data <= "000000";
--when "0100011001" => data <= "000000";
--when "0100011010" => data <= "000000";
--when "0100011011" => data <= "000000";
--when "0100011100" => data <= "000000";
--when "0101110100" => data <= "000000";
--when "0110000001" => data <= "000000";
--when "0110001000" => data <= "000000";
--when "0110001001" => data <= "000000";
		--when others => data <= "111111";
--end case;
--end process;
--end;











