library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity GameOverROM is
port(
	Xin : in unsigned(8 downto 0);
	Yin : in unsigned(8 downto 0);
data : out std_logic_vector(5 downto 0)
);
end GameOverROM;


architecture synth of GameOverROM is

signal addy : unsigned(17 downto 0);

begin

addy <= Yin & Xin;

process(addy) begin
	case addy is
when "000000000000000001" => data <= "000000";
when "000000000000000010" => data <= "000000";
when "000000000000000011" => data <= "000000";
when "000000000000000100" => data <= "000000";
when "000000000000001001" => data <= "000000";
when "000000000000001101" => data <= "000000";
when "000000000000001110" => data <= "000000";
when "000000000000001111" => data <= "000000";
when "000000000000010000" => data <= "000000";
when "000000000000010001" => data <= "000000";
when "000000000000010011" => data <= "000000";
when "000000000000010100" => data <= "000000";
when "000000000000010101" => data <= "000000";
when "000000000000010110" => data <= "000000";
when "000000000000100000" => data <= "000000";
when "000000000000100001" => data <= "000000";
when "000000000000100010" => data <= "000000";
when "000000000000100110" => data <= "000000";
when "000000000000101010" => data <= "000000";
when "000000000000101100" => data <= "000000";
when "000000000000101101" => data <= "000000";
when "000000000000101110" => data <= "000000";
when "000000000000101111" => data <= "000000";
when "000000000000110001" => data <= "000000";
when "000000000000110010" => data <= "000000";
when "000000000000110011" => data <= "000000";
when "000000000000110100" => data <= "000000";
when "000000001000000000" => data <= "000000";
when "000000001000000001" => data <= "000000";
when "000000001000001000" => data <= "000000";
when "000000001000001001" => data <= "000000";
when "000000001000001010" => data <= "000000";
when "000000001000001101" => data <= "000000";
when "000000001000001111" => data <= "000000";
when "000000001000010001" => data <= "000000";
when "000000001000010011" => data <= "000000";
when "000000001000011111" => data <= "000000";
when "000000001000100011" => data <= "000000";
when "000000001000100110" => data <= "000000";
when "000000001000101010" => data <= "000000";
when "000000001000101100" => data <= "000000";
when "000000001000110001" => data <= "000000";
when "000000001000110100" => data <= "000000";
when "000000010000000000" => data <= "000000";
when "000000010000001000" => data <= "000000";
when "000000010000001010" => data <= "000000";
when "000000010000001101" => data <= "000000";
when "000000010000001111" => data <= "000000";
when "000000010000010001" => data <= "000000";
when "000000010000010011" => data <= "000000";
when "000000010000011110" => data <= "000000";
when "000000010000100100" => data <= "000000";
when "000000010000100110" => data <= "000000";
when "000000010000101010" => data <= "000000";
when "000000010000101100" => data <= "000000";
when "000000010000110001" => data <= "000000";
when "000000010000110100" => data <= "000000";
when "000000011000000000" => data <= "000000";
when "000000011000000010" => data <= "000000";
when "000000011000000011" => data <= "000000";
when "000000011000000100" => data <= "000000";
when "000000011000000101" => data <= "000000";
when "000000011000000111" => data <= "000000";
when "000000011000001000" => data <= "000000";
when "000000011000001001" => data <= "000000";
when "000000011000001010" => data <= "000000";
when "000000011000001011" => data <= "000000";
when "000000011000001101" => data <= "000000";
when "000000011000001111" => data <= "000000";
when "000000011000010001" => data <= "000000";
when "000000011000010011" => data <= "000000";
when "000000011000010100" => data <= "000000";
when "000000011000010101" => data <= "000000";
when "000000011000010110" => data <= "000000";
when "000000011000011110" => data <= "000000";
when "000000011000100100" => data <= "000000";
when "000000011000100111" => data <= "000000";
when "000000011000101001" => data <= "000000";
when "000000011000101100" => data <= "000000";
when "000000011000101101" => data <= "000000";
when "000000011000101110" => data <= "000000";
when "000000011000101111" => data <= "000000";
when "000000011000110001" => data <= "000000";
when "000000011000110010" => data <= "000000";
when "000000011000110011" => data <= "000000";
when "000000011000110100" => data <= "000000";
when "000000100000000000" => data <= "000000";
when "000000100000000100" => data <= "000000";
when "000000100000000111" => data <= "000000";
when "000000100000001011" => data <= "000000";
when "000000100000001101" => data <= "000000";
when "000000100000010001" => data <= "000000";
when "000000100000010011" => data <= "000000";
when "000000100000011110" => data <= "000000";
when "000000100000100100" => data <= "000000";
when "000000100000100111" => data <= "000000";
when "000000100000101001" => data <= "000000";
when "000000100000101100" => data <= "000000";
when "000000100000110001" => data <= "000000";
when "000000100000110011" => data <= "000000";
when "000000101000000000" => data <= "000000";
when "000000101000000001" => data <= "000000";
when "000000101000000100" => data <= "000000";
when "000000101000000111" => data <= "000000";
when "000000101000001011" => data <= "000000";
when "000000101000001101" => data <= "000000";
when "000000101000010001" => data <= "000000";
when "000000101000010011" => data <= "000000";
when "000000101000011111" => data <= "000000";
when "000000101000100011" => data <= "000000";
when "000000101000100111" => data <= "000000";
when "000000101000101000" => data <= "000000";
when "000000101000101001" => data <= "000000";
when "000000101000101100" => data <= "000000";
when "000000101000110001" => data <= "000000";
when "000000101000110100" => data <= "000000";
when "000000110000000001" => data <= "000000";
when "000000110000000010" => data <= "000000";
when "000000110000000011" => data <= "000000";
when "000000110000000100" => data <= "000000";
when "000000110000000111" => data <= "000000";
when "000000110000001011" => data <= "000000";
when "000000110000001101" => data <= "000000";
when "000000110000010001" => data <= "000000";
when "000000110000010011" => data <= "000000";
when "000000110000010100" => data <= "000000";
when "000000110000010101" => data <= "000000";
when "000000110000010110" => data <= "000000";
when "000000110000100000" => data <= "000000";
when "000000110000100001" => data <= "000000";
when "000000110000100010" => data <= "000000";
when "000000110000101000" => data <= "000000";
when "000000110000101100" => data <= "000000";
when "000000110000101101" => data <= "000000";
when "000000110000101110" => data <= "000000";
when "000000110000101111" => data <= "000000";
when "000000110000110001" => data <= "000000";
when "000000110000110100" => data <= "000000";
when "000001100000010101" => data <= "000000";
when "000001100000010110" => data <= "000000";
when "000001100000010111" => data <= "000000";
when "000001100000011000" => data <= "000000";
when "000001100000011001" => data <= "000000";
when "000001100000011010" => data <= "000000";
when "000001100000011011" => data <= "000000";
when "000001100000011100" => data <= "000000";
when "000001100000011101" => data <= "000000";
when "000001100000011110" => data <= "000000";
when "000001100000011111" => data <= "000000";
when "000001100000100000" => data <= "000000";
when "000001100000100001" => data <= "000000";
when "000001101000010101" => data <= "000000";
when "000001101000010110" => data <= "000000";
when "000001101000010111" => data <= "000000";
when "000001101000011000" => data <= "000000";
when "000001101000011010" => data <= "000000";
when "000001101000011011" => data <= "000000";
when "000001101000011100" => data <= "000000";
when "000001101000011101" => data <= "000000";
when "000001101000011110" => data <= "000000";
when "000001101000011111" => data <= "000000";
when "000001101000100000" => data <= "000000";
when "000001101000100001" => data <= "000000";
when "000001110000010101" => data <= "000000";
when "000001110000010110" => data <= "000000";
when "000001110000010111" => data <= "000000";
when "000001110000011000" => data <= "000000";
when "000001110000011011" => data <= "000000";
when "000001110000011100" => data <= "000000";
when "000001110000011101" => data <= "000000";
when "000001110000011110" => data <= "000000";
when "000001110000011111" => data <= "000000";
when "000001110000100000" => data <= "000000";
when "000001110000100001" => data <= "000000";
when "000001111000010101" => data <= "000000";
when "000001111000010110" => data <= "000000";
when "000001111000011100" => data <= "000000";
when "000001111000100000" => data <= "000000";
when "000001111000100001" => data <= "000000";
when "000010000000010101" => data <= "000000";
when "000010000000010110" => data <= "000000";
when "000010000000011000" => data <= "000000";
when "000010000000011011" => data <= "000000";
when "000010000000011100" => data <= "000000";
when "000010000000011101" => data <= "000000";
when "000010000000011110" => data <= "000000";
when "000010000000100000" => data <= "000000";
when "000010000000100001" => data <= "000000";
when "000010001000010101" => data <= "000000";
when "000010001000010110" => data <= "000000";
when "000010001000011000" => data <= "000000";
when "000010001000011010" => data <= "000000";
when "000010001000011011" => data <= "000000";
when "000010001000011100" => data <= "000000";
when "000010001000011101" => data <= "000000";
when "000010001000011110" => data <= "000000";
when "000010001000100000" => data <= "000000";
when "000010001000100001" => data <= "000000";
when "000010010000010101" => data <= "000000";
when "000010010000010110" => data <= "000000";
when "000010010000011000" => data <= "000000";
when "000010010000011001" => data <= "000000";
when "000010010000011010" => data <= "000000";
when "000010010000011011" => data <= "000000";
when "000010010000011100" => data <= "000000";
when "000010010000011101" => data <= "000000";
when "000010010000011110" => data <= "000000";
when "000010010000100000" => data <= "000000";
when "000010010000100001" => data <= "000000";
when "000010011000010101" => data <= "000000";
when "000010011000010110" => data <= "000000";
when "000010011000011000" => data <= "000000";
when "000010011000011001" => data <= "000000";
when "000010011000011010" => data <= "000000";
when "000010011000011011" => data <= "000000";
when "000010011000011100" => data <= "000000";
when "000010011000011101" => data <= "000000";
when "000010011000011110" => data <= "000000";
when "000010011000100000" => data <= "000000";
when "000010011000100001" => data <= "000000";
when "000010100000010101" => data <= "000000";
when "000010100000010110" => data <= "000000";
when "000010100000011000" => data <= "000000";
when "000010100000011001" => data <= "000000";
when "000010100000011010" => data <= "000000";
when "000010100000011011" => data <= "000000";
when "000010100000011100" => data <= "000000";
when "000010100000011101" => data <= "000000";
when "000010100000011110" => data <= "000000";
when "000010100000100000" => data <= "000000";
when "000010100000100001" => data <= "000000";
when "000010101000010101" => data <= "000000";
when "000010101000010110" => data <= "000000";
when "000010101000100000" => data <= "000000";
when "000010101000100001" => data <= "000000";
when "000010110000010101" => data <= "000000";
when "000010110000010110" => data <= "000000";
when "000010110000010111" => data <= "000000";
when "000010110000011000" => data <= "000000";
when "000010110000011001" => data <= "000000";
when "000010110000011010" => data <= "000000";
when "000010110000011011" => data <= "000000";
when "000010110000011100" => data <= "000000";
when "000010110000011101" => data <= "000000";
when "000010110000011110" => data <= "000000";
when "000010110000011111" => data <= "000000";
when "000010110000100000" => data <= "000000";
when "000010110000100001" => data <= "000000";
when "000010111000010101" => data <= "000000";
when "000010111000010110" => data <= "000000";
when "000010111000010111" => data <= "000000";
when "000010111000011000" => data <= "000000";
when "000010111000011001" => data <= "000000";
when "000010111000011010" => data <= "000000";
when "000010111000011011" => data <= "000000";
when "000010111000011100" => data <= "000000";
when "000010111000011101" => data <= "000000";
when "000010111000011110" => data <= "000000";
when "000010111000011111" => data <= "000000";
when "000010111000100000" => data <= "000000";
when "000010111000100001" => data <= "000000";

when others => data <= "111111";

end case;
end process;
end;
