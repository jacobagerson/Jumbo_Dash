--library IEEE;
--use IEEE.std_logic_1164.all;
--use IEEE.numeric_std.all;


--entity ground1ROM is
--port(
	--Xin : in unsigned(4 downto 0);
	--Yin : in unsigned(4 downto 0);
--data : out std_logic_vector(5 downto 0)
--);
--end entity;


--architecture synth of ground1ROM is


--Signal addy : unsigned(9 downto 0);


--Begin


--addy <= Yin & Xin;


--process(addy) begin
	--case addy is
		--when "0001100000" => data <= "000000";
--when "0001100001" => data <= "000000";
--when "0001100010" => data <= "000000";
--when "0001100011" => data <= "000000";
--when "0001100100" => data <= "000000";
--when "0001100101" => data <= "000000";
--when "0001100110" => data <= "000000";
--when "0001100111" => data <= "000000";
--when "0001101000" => data <= "000000";
--when "0001101001" => data <= "000000";
--when "0001101010" => data <= "000000";
--when "0001101011" => data <= "000000";
--when "0001101100" => data <= "000000";
--when "0001101101" => data <= "000000";
--when "0001101110" => data <= "000000";
--when "0001101111" => data <= "000000";
--when "0001110000" => data <= "000000";
--when "0001110001" => data <= "000000";
--when "0001110010" => data <= "000000";
--when "0001110011" => data <= "000000";
--when "0001110100" => data <= "000000";
--when "0001110101" => data <= "000000";
--when "0001110110" => data <= "000000";
--when "0001110111" => data <= "000000";
--when "0001111000" => data <= "000000";
--when "0001111001" => data <= "000000";
--when "0001111010" => data <= "000000";
--when "0001111011" => data <= "000000";
--when "0001111100" => data <= "000000";
--when "0001111101" => data <= "000000";
--when "0001111110" => data <= "000000";
--when "0011000101" => data <= "000000";
--when "0011000110" => data <= "000000";
--when "0011000111" => data <= "000000";
--when "0011011010" => data <= "000000";
--when "0011011011" => data <= "000000";
--when "0100001110" => data <= "000000";
--when "0111001011" => data <= "000000";
--when "0111001100" => data <= "000000";
		--when others => data <= "111111";
--end case;
--end process;
--end;











