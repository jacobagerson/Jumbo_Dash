library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity biggroundROM is
port(
Xin : in unsigned(8 downto 0);
Yin : in unsigned(8 downto 0);
data : out std_logic_vector(5 downto 0)
);
end entity;


architecture synth of biggroundROM is


Signal addy : unsigned(17 downto 0);


begin


addy <= Yin & Xin;


process(addy) begin
	case addy is
when "000000000010100111" => data <= "000000";
when "000000000010101000" => data <= "000000";
when "000000000010101001" => data <= "000000";
when "000000000010101010" => data <= "000000";
when "000000000010101011" => data <= "000000";
when "000000000010101100" => data <= "000000";
when "000000000010101101" => data <= "000000";
when "000000000010101110" => data <= "000000";
when "000000000010101111" => data <= "000000";
when "000000000010110000" => data <= "000000";
when "000000000010110001" => data <= "000000";
when "000000001010100110" => data <= "000000";
when "000000001010100111" => data <= "000000";
when "000000001010110001" => data <= "000000";
when "000000001010110010" => data <= "000000";
when "000000010010100101" => data <= "000000";
when "000000010010100110" => data <= "000000";
when "000000010010110010" => data <= "000000";
when "000000010010110011" => data <= "000000";
when "000000011010100100" => data <= "000000";
when "000000011010100101" => data <= "000000";
when "000000011010110011" => data <= "000000";
when "000000011100100111" => data <= "000000";
when "000000011100101000" => data <= "000000";
when "000000011100101001" => data <= "000000";
when "000000011100101010" => data <= "000000";
when "000000100001011101" => data <= "000000";
when "000000100001011110" => data <= "000000";
when "000000100001011111" => data <= "000000";
when "000000100001100000" => data <= "000000";
when "000000100001100001" => data <= "000000";
when "000000100001100010" => data <= "000000";
when "000000100001100011" => data <= "000000";
when "000000100001100100" => data <= "000000";
when "000000100001100101" => data <= "000000";
when "000000100001100110" => data <= "000000";
when "000000100010100001" => data <= "000000";
when "000000100010100010" => data <= "000000";
when "000000100010100011" => data <= "000000";
when "000000100010100100" => data <= "000000";
when "000000100010110011" => data <= "000000";
when "000000100010110100" => data <= "000000";
when "000000100010110101" => data <= "000000";
when "000000100010110110" => data <= "000000";
when "000000100100100110" => data <= "000000";
when "000000100100100111" => data <= "000000";
when "000000100100101010" => data <= "000000";
when "000000100100101011" => data <= "000000";
when "000000101001011100" => data <= "000000";
when "000000101001011101" => data <= "000000";
when "000000101001100110" => data <= "000000";
when "000000101001100111" => data <= "000000";
when "000000101010100000" => data <= "000000";
when "000000101010100001" => data <= "000000";
when "000000101010110110" => data <= "000000";
when "000000101010110111" => data <= "000000";
when "000000101100100000" => data <= "000000";
when "000000101100100001" => data <= "000000";
when "000000101100100010" => data <= "000000";
when "000000101100100011" => data <= "000000";
when "000000101100100100" => data <= "000000";
when "000000101100100101" => data <= "000000";
when "000000101100100110" => data <= "000000";
when "000000101100101011" => data <= "000000";
when "000000101100101100" => data <= "000000";
when "000000101100101101" => data <= "000000";
when "000000101100101110" => data <= "000000";
when "000000110000000000" => data <= "000000";
when "000000110000000001" => data <= "000000";
when "000000110000000010" => data <= "000000";
when "000000110000000011" => data <= "000000";
when "000000110000000100" => data <= "000000";
when "000000110000000101" => data <= "000000";
when "000000110000000110" => data <= "000000";
when "000000110000000111" => data <= "000000";
when "000000110000001000" => data <= "000000";
when "000000110000001001" => data <= "000000";
when "000000110000001010" => data <= "000000";
when "000000110000001011" => data <= "000000";
when "000000110000001100" => data <= "000000";
when "000000110000001101" => data <= "000000";
when "000000110000001110" => data <= "000000";
when "000000110000001111" => data <= "000000";
when "000000110000010000" => data <= "000000";
when "000000110000010001" => data <= "000000";
when "000000110000010010" => data <= "000000";
when "000000110000010011" => data <= "000000";
when "000000110000010100" => data <= "000000";
when "000000110000010101" => data <= "000000";
when "000000110000010110" => data <= "000000";
when "000000110000010111" => data <= "000000";
when "000000110000011000" => data <= "000000";
when "000000110000011001" => data <= "000000";
when "000000110000011010" => data <= "000000";
when "000000110000011011" => data <= "000000";
when "000000110000011100" => data <= "000000";
when "000000110000011101" => data <= "000000";
when "000000110000011110" => data <= "000000";
when "000000110000011111" => data <= "000000";
when "000000110000100000" => data <= "000000";
when "000000110000100001" => data <= "000000";
when "000000110000100010" => data <= "000000";
when "000000110000100011" => data <= "000000";
when "000000110000100100" => data <= "000000";
when "000000110000100101" => data <= "000000";
when "000000110000100110" => data <= "000000";
when "000000110000100111" => data <= "000000";
when "000000110000101000" => data <= "000000";
when "000000110000101001" => data <= "000000";
when "000000110000101010" => data <= "000000";
when "000000110000101011" => data <= "000000";
when "000000110000101100" => data <= "000000";
when "000000110000101101" => data <= "000000";
when "000000110000101110" => data <= "000000";
when "000000110000101111" => data <= "000000";
when "000000110000110000" => data <= "000000";
when "000000110000110001" => data <= "000000";
when "000000110000110010" => data <= "000000";
when "000000110000110011" => data <= "000000";
when "000000110000110100" => data <= "000000";
when "000000110000110101" => data <= "000000";
when "000000110000110110" => data <= "000000";
when "000000110000110111" => data <= "000000";
when "000000110000111000" => data <= "000000";
when "000000110000111001" => data <= "000000";
when "000000110000111010" => data <= "000000";
when "000000110000111011" => data <= "000000";
when "000000110000111100" => data <= "000000";
when "000000110000111101" => data <= "000000";
when "000000110000111110" => data <= "000000";
when "000000110000111111" => data <= "000000";
when "000000110001000000" => data <= "000000";
when "000000110001000001" => data <= "000000";
when "000000110001000010" => data <= "000000";
when "000000110001000011" => data <= "000000";
when "000000110001000100" => data <= "000000";
when "000000110001000101" => data <= "000000";
when "000000110001000110" => data <= "000000";
when "000000110001000111" => data <= "000000";
when "000000110001001000" => data <= "000000";
when "000000110001001001" => data <= "000000";
when "000000110001001010" => data <= "000000";
when "000000110001001011" => data <= "000000";
when "000000110001001100" => data <= "000000";
when "000000110001001101" => data <= "000000";
when "000000110001001110" => data <= "000000";
when "000000110001001111" => data <= "000000";
when "000000110001011011" => data <= "000000";
when "000000110001011100" => data <= "000000";
when "000000110001100111" => data <= "000000";
when "000000110001101000" => data <= "000000";
when "000000110001101001" => data <= "000000";
when "000000110001101010" => data <= "000000";
when "000000110001101011" => data <= "000000";
when "000000110001101100" => data <= "000000";
when "000000110001101101" => data <= "000000";
when "000000110001101110" => data <= "000000";
when "000000110001101111" => data <= "000000";
when "000000110001110000" => data <= "000000";
when "000000110001110001" => data <= "000000";
when "000000110001110010" => data <= "000000";
when "000000110001110011" => data <= "000000";
when "000000110001110100" => data <= "000000";
when "000000110001110101" => data <= "000000";
when "000000110001110110" => data <= "000000";
when "000000110001110111" => data <= "000000";
when "000000110001111000" => data <= "000000";
when "000000110001111001" => data <= "000000";
when "000000110001111010" => data <= "000000";
when "000000110001111011" => data <= "000000";
when "000000110001111100" => data <= "000000";
when "000000110001111101" => data <= "000000";
when "000000110001111110" => data <= "000000";
when "000000110001111111" => data <= "000000";
when "000000110010000000" => data <= "000000";
when "000000110010000001" => data <= "000000";
when "000000110010000010" => data <= "000000";
when "000000110010000011" => data <= "000000";
when "000000110010000100" => data <= "000000";
when "000000110010000101" => data <= "000000";
when "000000110010000110" => data <= "000000";
when "000000110010000111" => data <= "000000";
when "000000110010001000" => data <= "000000";
when "000000110010001001" => data <= "000000";
when "000000110010001010" => data <= "000000";
when "000000110010001011" => data <= "000000";
when "000000110010001100" => data <= "000000";
when "000000110010001101" => data <= "000000";
when "000000110010001110" => data <= "000000";
when "000000110010001111" => data <= "000000";
when "000000110010010000" => data <= "000000";
when "000000110010010001" => data <= "000000";
when "000000110010010010" => data <= "000000";
when "000000110010010011" => data <= "000000";
when "000000110010010100" => data <= "000000";
when "000000110010010101" => data <= "000000";
when "000000110010010110" => data <= "000000";
when "000000110010010111" => data <= "000000";
when "000000110010011000" => data <= "000000";
when "000000110010011001" => data <= "000000";
when "000000110010011010" => data <= "000000";
when "000000110010011011" => data <= "000000";
when "000000110010011100" => data <= "000000";
when "000000110010011101" => data <= "000000";
when "000000110010011110" => data <= "000000";
when "000000110010011111" => data <= "000000";
when "000000110010100000" => data <= "000000";
when "000000110010110111" => data <= "000000";
when "000000110010111000" => data <= "000000";
when "000000110010111001" => data <= "000000";
when "000000110010111010" => data <= "000000";
when "000000110010111011" => data <= "000000";
when "000000110010111100" => data <= "000000";
when "000000110010111101" => data <= "000000";
when "000000110010111110" => data <= "000000";
when "000000110010111111" => data <= "000000";
when "000000110011000000" => data <= "000000";
when "000000110011000001" => data <= "000000";
when "000000110011000010" => data <= "000000";
when "000000110011000011" => data <= "000000";
when "000000110011000100" => data <= "000000";
when "000000110011000101" => data <= "000000";
when "000000110011000110" => data <= "000000";
when "000000110011000111" => data <= "000000";
when "000000110011001000" => data <= "000000";
when "000000110011001001" => data <= "000000";
when "000000110011001010" => data <= "000000";
when "000000110011001011" => data <= "000000";
when "000000110011001100" => data <= "000000";
when "000000110011001101" => data <= "000000";
when "000000110011001110" => data <= "000000";
when "000000110011001111" => data <= "000000";
when "000000110011010000" => data <= "000000";
when "000000110011010001" => data <= "000000";
when "000000110011010010" => data <= "000000";
when "000000110011010011" => data <= "000000";
when "000000110011010100" => data <= "000000";
when "000000110011010101" => data <= "000000";
when "000000110011010110" => data <= "000000";
when "000000110011010111" => data <= "000000";
when "000000110011011000" => data <= "000000";
when "000000110011011001" => data <= "000000";
when "000000110011011010" => data <= "000000";
when "000000110011011011" => data <= "000000";
when "000000110011011100" => data <= "000000";
when "000000110011011101" => data <= "000000";
when "000000110011011110" => data <= "000000";
when "000000110011011111" => data <= "000000";
when "000000110011100000" => data <= "000000";
when "000000110011100001" => data <= "000000";
when "000000110011100010" => data <= "000000";
when "000000110011100011" => data <= "000000";
when "000000110011100100" => data <= "000000";
when "000000110011100101" => data <= "000000";
when "000000110011100110" => data <= "000000";
when "000000110011100111" => data <= "000000";
when "000000110011101000" => data <= "000000";
when "000000110011101001" => data <= "000000";
when "000000110011101010" => data <= "000000";
when "000000110011101011" => data <= "000000";
when "000000110011101100" => data <= "000000";
when "000000110011101101" => data <= "000000";
when "000000110011101110" => data <= "000000";
when "000000110011101111" => data <= "000000";
when "000000110011110000" => data <= "000000";
when "000000110011110001" => data <= "000000";
when "000000110011110010" => data <= "000000";
when "000000110011110011" => data <= "000000";
when "000000110011110100" => data <= "000000";
when "000000110011110101" => data <= "000000";
when "000000110100000010" => data <= "000000";
when "000000110100000011" => data <= "000000";
when "000000110100000100" => data <= "000000";
when "000000110100000101" => data <= "000000";
when "000000110100000110" => data <= "000000";
when "000000110100000111" => data <= "000000";
when "000000110100001000" => data <= "000000";
when "000000110100001001" => data <= "000000";
when "000000110100001010" => data <= "000000";
when "000000110100001011" => data <= "000000";
when "000000110100001100" => data <= "000000";
when "000000110100001101" => data <= "000000";
when "000000110100001110" => data <= "000000";
when "000000110100001111" => data <= "000000";
when "000000110100010000" => data <= "000000";
when "000000110100010001" => data <= "000000";
when "000000110100010010" => data <= "000000";
when "000000110100010011" => data <= "000000";
when "000000110100010100" => data <= "000000";
when "000000110100010101" => data <= "000000";
when "000000110100010110" => data <= "000000";
when "000000110100010111" => data <= "000000";
when "000000110100011000" => data <= "000000";
when "000000110100011001" => data <= "000000";
when "000000110100011010" => data <= "000000";
when "000000110100011011" => data <= "000000";
when "000000110100011100" => data <= "000000";
when "000000110100011101" => data <= "000000";
when "000000110100011110" => data <= "000000";
when "000000110100011111" => data <= "000000";
when "000000110100100000" => data <= "000000";
when "000000110100101110" => data <= "000000";
when "000000110100101111" => data <= "000000";
when "000000110100110000" => data <= "000000";
when "000000110100110001" => data <= "000000";
when "000000110100110010" => data <= "000000";
when "000000110100110011" => data <= "000000";
when "000000110100110100" => data <= "000000";
when "000000110100110101" => data <= "000000";
when "000000110100110110" => data <= "000000";
when "000000110100110111" => data <= "000000";
when "000000110100111000" => data <= "000000";
when "000000110100111001" => data <= "000000";
when "000000110100111010" => data <= "000000";
when "000000110100111011" => data <= "000000";
when "000000110100111100" => data <= "000000";
when "000000110100111101" => data <= "000000";
when "000000110100111110" => data <= "000000";
when "000000110100111111" => data <= "000000";
when "000000111001001111" => data <= "000000";
when "000000111001011010" => data <= "000000";
when "000000111001011011" => data <= "000000";
when "000000111011110101" => data <= "000000";
when "000000111011110110" => data <= "000000";
when "000000111100000001" => data <= "000000";
when "000000111100000010" => data <= "000000";
when "000001000001001111" => data <= "000000";
when "000001000001010000" => data <= "000000";
when "000001000001010001" => data <= "000000";
when "000001000001010010" => data <= "000000";
when "000001000001010011" => data <= "000000";
when "000001000001010100" => data <= "000000";
when "000001000001010101" => data <= "000000";
when "000001000001010110" => data <= "000000";
when "000001000001010111" => data <= "000000";
when "000001000001011000" => data <= "000000";
when "000001000001011001" => data <= "000000";
when "000001000001011010" => data <= "000000";
when "000001000011110110" => data <= "000000";
when "000001000011110111" => data <= "000000";
when "000001000011111000" => data <= "000000";
when "000001000011111001" => data <= "000000";
when "000001000011111010" => data <= "000000";
when "000001000011111011" => data <= "000000";
when "000001000011111100" => data <= "000000";
when "000001000011111101" => data <= "000000";
when "000001000011111110" => data <= "000000";
when "000001000011111111" => data <= "000000";
when "000001000100000000" => data <= "000000";
when "000001000100000001" => data <= "000000";
when "000001101000001010" => data <= "000000";
when "000001101000001011" => data <= "000000";
when "000001101000001100" => data <= "000000";
when "000001101000001101" => data <= "000000";
when "000001101000001110" => data <= "000000";
when "000001101000110100" => data <= "000000";
when "000001101000110101" => data <= "000000";
when "000001101000110110" => data <= "000000";
when "000001101000110111" => data <= "000000";
when "000001101001110010" => data <= "000000";
when "000001101001110011" => data <= "000000";
when "000001101001110100" => data <= "000000";
when "000001101001110101" => data <= "000000";
when "000001101100101001" => data <= "000000";
when "000001101100101010" => data <= "000000";
when "000001111010100100" => data <= "000000";
when "000001111010100101" => data <= "000000";
when "000010000011011000" => data <= "000000";
when "000010000011011001" => data <= "000000";
when "000010001000011100" => data <= "000000";
when "000010001010000010" => data <= "000000";
when "000010001010000011" => data <= "000000";
when "000010010100011000" => data <= "000000";
when "000010010100011001" => data <= "000000";
when "000010010100011010" => data <= "000000";
when "000010010100011011" => data <= "000000";
when "000010011001001100" => data <= "000000";
when "000010011001001101" => data <= "000000";
when "000010011001001110" => data <= "000000";
when "000010011001001111" => data <= "000000";
when "000010011001010000" => data <= "000000";
when "000010011001010001" => data <= "000000";
when "000010011010111010" => data <= "000000";
when "000010011010111011" => data <= "000000";
when "000010011010111100" => data <= "000000";
when "000010011010111101" => data <= "000000";
when "000010011011110010" => data <= "000000";
when "000010011011110011" => data <= "000000";
when "000010101001100000" => data <= "000000";
when "000010101001100001" => data <= "000000";
when "000010111010011010" => data <= "000000";
when "000010111100110010" => data <= "000000";
when "000010111100110011" => data <= "000000";
when "000010111100110100" => data <= "000000";
when "000010111100110101" => data <= "000000";
when "000011001011000010" => data <= "000000";
when "000011001011000011" => data <= "000000";
when "000011001011000100" => data <= "000000";
when "000011011011101100" => data <= "000000";
when "000011011011101101" => data <= "000000";
when "000011011011101110" => data <= "000000";
when "000011011011101111" => data <= "000000";
when "000011011011110000" => data <= "000000";
when "000011011011110001" => data <= "000000";
when "000011101000010110" => data <= "000000";
when "000011101000010111" => data <= "000000";
when "000011101000011000" => data <= "000000";
when "000011101000011001" => data <= "000000";
when "000011101100010110" => data <= "000000";








		when others => data <= "111111";
end case;
end process;
end;

